`timescale 1ns / 1ps

module EXU32 #(  //EXecution Unit
    INST_MAX = 32,
    WIDTH    = 32
) ();
endmodule
