`timescale 1ns / 1ps

module Multiplier #(  //快速乘法器
    WIDTH = 32
) (
    input  [  WIDTH-1:0] in1,
    input  [  WIDTH-1:0] in2,
    output [WIDTH*2-1:0] out
);

endmodule
